LastName ! FirstName ! Gender ! FavoriteColor ! DateOfBirth
Einstein ! Albert ! Male ! Green ! 03/14/1879
Darwin ! Charles ! Male ! Blue ! 02/12/1809
Curie ! Marie ! Female ! Yellow ! 11/07/1867
Lovelace ! Ada ! Female ! Purple ! 12/10/1815
Turing ! Alan ! Male ! Red ! 06/03/1912
