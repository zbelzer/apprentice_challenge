LastName ! FirstName ! Gender ! FavoriteColor ! DateOfBirth
Einstein ! Albert ! Male ! Green ! 1879-03-14
Darwin ! Charles ! Male ! Blue ! 1809-02-12
Curie ! Marie ! Female ! Yellow ! 1867-11-07
Lovelace ! Ada ! Female ! Purple ! 1815-12-10
Turing ! Alan ! Male ! Red ! 1912-06-03
